library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity DF is 
port(
			reset		: in std_logic;
			mode		: in std_logic;
			increase : in std_logic;
			decrease : in std_logic;
			clock_400: in std_logic


);
end entity DF;

architecture rtl of DF is 
begin

end architecture rtl;