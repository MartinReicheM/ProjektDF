library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity DigitalFilter is 
port(
		input : in std_logic
);
end entity;

architecture rtl of DigitalFilter is 

begin 

end architecture rtl;
